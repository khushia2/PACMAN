module characters_rom (
    input [5:0] addr,
    output [15:0] data
);

parameter ADDR_WIDTH = 6;
parameter DATA_WIDTH =  16;

logic [ADDR_WIDTH-1:0] addr_reg;

parameter [0:47][DATA_WIDTH-1:0] ROM = {
    //GHOST
    16'b0000000000000000,
    16'b0000111111110000,
    16'b0111111111111110,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111000111100011,
    16'b1111000111100011,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1101111001111011,
    16'b1000110000110001,
    //PACMAN - OPEN
    16'b0000000000000000,
    16'b0000011111100000,
    16'b0001111111111000,
    16'b0011111100011100,
    16'b0111111100011110,
    16'b1111111111111110,
    16'b1111111111100000,
    16'b1111111000000000,
    16'b1111111000000000,
    16'b1111111111100000,
    16'b1111111111111110,
    16'b0111111111111110,
    16'b0011111111111100,
    16'b0001111111111000,
    16'b0000011111100000,
    16'b0000000000000000,
    //PACMAN - CLOSED
    16'b0000000000000000,
    16'b0000011111100000,
    16'b0001111111111000,
    16'b0011111100011100,
    16'b0111111100011110,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b1111111111111111,
    16'b0111111111111110,
    16'b0011111111111100,
    16'b0001111111111000,
    16'b0000011111100000,
    16'b0000000000000000,
};

assign data = ROM[addr];

endmodule