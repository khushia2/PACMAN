module maze_array_rom (
    input [8:0] addr,
    output [0:639] data
);

parameter ADDR_WIDTH = 9;
parameter DATA_WIDTH = 640;

parameter logic [0:DATA_WIDTH-1] ROM [0:479] = '{
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    -640'd1,
    -640'd1,
    -640'd1,
    -640'd1,
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -91'd1, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, -119'd1, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -91'd1, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, -119'd1, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -91'd1, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, -119'd1, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -91'd1, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, -119'd1, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b0, 18'b0, 75'b0, 18'b0, 91'b0, 18'b0, 4'b1111, 72'b0, 4'b1111, 18'b0, 119'b0, 18'b0, 75'b0, 18'b0, 4'b0, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -91'd1, 18'b0, -80'd1, 18'b0, -119'd1, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -91'd1, 18'b0, -80'd1, 18'b0, -119'd1, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -91'd1, 18'b0, -80'd1, 18'b0, -119'd1, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -91'd1, 18'b0, -80'd1, 18'b0, -119'd1, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b0, 362'b0, 4'b0, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 362'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -53'd1, 18'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, 4'b1111, 89'b0, 4'b1111, 362'b0, 4'b1111, 89'b0, 4'b1111, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -34'd1},
    {10'b0, 4'b1111, 18'b0, -75'd1, 18'b0, 4'b1111, 18'b0, -326'd1, 18'b0, 4'b1111, 18'b0, -75'd1, 18'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    {10'b0, 4'b1111, 111'b0, 4'b1111, 362'b0, 4'b1111, 111'b0, -34'd1},
    -640'd1,
    -640'd1,
    -640'd1,
    -640'd1,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0,
    640'b0
};

assign data = ROM[addr];

endmodule