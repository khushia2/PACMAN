module bigfont_rom (
    input [8:0]	addr,
	output [23:0]	data
);

parameter ADDR_WIDTH = 9;
parameter DATA_WIDTH =  24;

logic [ADDR_WIDTH-1:0] addr_reg;

parameter [0:319][DATA_WIDTH-1:0] ROM = {
    //P
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,   
    24'b111111111111111111000000,
    24'b111111111111111111000000,
    24'b111111111111111111000000, 
    24'b000111111000000111111000, 
    24'b000111111000000111111000, 
    24'b000111111000000111111000, 
    24'b000111111000000111111000, 
    24'b000111111000000111111000,
    24'b000111111000000111111000, 
    24'b000111111000000111111000, 
    24'b000111111000000111111000,
    24'b000111111000000111111000,   
    24'b000111111111111111000000, 
    24'b000111111111111111000000, 
    24'b000111111111111111000000, 
    24'b000111111000000000000000, 
    24'b000111111000000000000000, 
    24'b000111111000000000000000, 
    24'b000111111000000000000000,
    24'b000111111000000000000000, 
    24'b000111111000000000000000, 
    24'b000111111000000000000000, 
    24'b000111111000000000000000,
    24'b000111111000000000000000, 
    24'b000111111000000000000000, 
    24'b000111111000000000000000, 
    24'b000111111000000000000000, 
    24'b111111111111000000000000,
    24'b111111111111000000000000, 
    24'b111111111111000000000000,  
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    //A
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000111000000000000,
    24'b000000000111000000000000,
    24'b000000000111000000000000,
    24'b000000111111111000000000,
    24'b000000111111111000000000,
    24'b000000111111111000000000,
    24'b000111111000111111000000,
    24'b000111111000111111000000,
    24'b000111111000111111000000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111111111111111111000,
    24'b111111111111111111111000,
    24'b111111111111111111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b111111000000000111111000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    //C
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000111111111111000000,
    24'b000000111111111111000000,
    24'b000000111111111111000000,
    24'b000111111000000111111000,
    24'b000111111000000111111000,
    24'b000111111000000111111000,
    24'b111111000000000000111000,
    24'b111111000000000000111000,
    24'b111111000000000000111000,
    24'b111111000000000000000000,
    24'b111111000000000000000000,
    24'b111111000000000000000000,
    24'b111111000000000000000000,
    24'b111111000000000000000000,
    24'b111111000000000000000000,
    24'b111111000000000000000000,
    24'b111111000000000000000000,
    24'b111111000000000000000000,
    24'b111111000000000000000000,
    24'b111111000000000000000000,
    24'b111111000000000000000000,
    24'b111111000000000000111000,
    24'b111111000000000000111000,
    24'b111111000000000000111000,
    24'b000111111000000111111000,
    24'b000111111000000111111000,
    24'b000111111000000111111000,
    24'b000000111111111111000000,
    24'b000000111111111111000000,
    24'b000000111111111111000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    //M
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111111000000000000111111,
    24'b111111000000000000111111,
    24'b111111000000000000111111,
    24'b111111111000000111111111,
    24'b111111111000000111111111,
    24'b111111111000000111111111,
    24'b111111111111111111111111, 
    24'b111111111111111111111111,
    24'b111111111111111111111111, 
    24'b111111111111111111111111,
    24'b111111111111111111111111, 
    24'b111111111111111111111111, 
    24'b111111000111111000111111,
    24'b111111000111111000111111, 
    24'b111111000111111000111111,  
    24'b111111000000000000111111, 
    24'b111111000000000000111111,
    24'b111111000000000000111111, 
    24'b111111000000000000111111, 
    24'b111111000000000000111111,
    24'b111111000000000000111111, 
    24'b111111000000000000111111,
    24'b111111000000000000111111, 
    24'b111111000000000000111111, 
    24'b111111000000000000111111,
    24'b111111000000000000111111, 
    24'b111111000000000000111111,
    24'b111111000000000000111111, 
    24'b111111000000000000111111, 
    24'b111111000000000000111111, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    //N
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b111111000000000111111000, 
    24'b111111000000000111111000, 
    24'b111111000000000111111000, 
    24'b111111111000000111111000, 
    24'b111111111000000111111000, 
    24'b111111111000000111111000, 
    24'b111111111111000111111000, 
    24'b111111111111000111111000,
    24'b111111111111000111111000,
    24'b111111111111111111111000, 
    24'b111111111111111111111000, 
    24'b111111111111111111111000, 
    24'b111111000111111111111000, 
    24'b111111000111111111111000, 
    24'b111111000111111111111000, 
    24'b111111000000111111111000, 
    24'b111111000000111111111000,
    24'b111111000000111111111000,
    24'b111111000000000111111000, 
    24'b111111000000000111111000, 
    24'b111111000000000111111000, 
    24'b111111000000000111111000,
    24'b111111000000000111111000, 
    24'b111111000000000111111000, 
    24'b111111000000000111111000, 
    24'b111111000000000111111000, 
    24'b111111000000000111111000, 
    24'b111111000000000111111000, 
    24'b111111000000000111111000, 
    24'b111111000000000111111000,  
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000,
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000, 
    24'b000000000000000000000000 
}; 

assign data = ROM[addr];

endmodule