module special_walls_2_rom (
    input [7:0] addr,
    output [3:0] data
);

parameter ADDR_WIDTH = 8;
parameter DATA_WIDTH = 4;

logic [ADDR_WIDTH-1:0] addr_reg;

parameter [0:166][DATA_WIDTH-1:0] ROM = {
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
};

assign data = ROM[addr];

endmodule