module special_walls_1_rom (
    input [4:0] addr,
    output [79:0] data
);

parameter ADDR_WIDTH = 5;
parameter DATA_WIDTH = 80;

logic [ADDR_WIDTH-1:0] addr_reg;

parameter [0:25][DATA_WIDTH-1:0] ROM = {
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111,
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111,
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111,
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111,
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111,
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111,
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111, 
    80'b11110000000000000000000000000000000000000000000000000000000000000000000000001111,
    -80'd1,
    -80'd1,
    -80'd1,
    -80'd1
};

assign data = ROM[addr];

endmodule