module special_walls_5_rom (
    input [9:0] addr,
    output [74:0] data
);

parameter ADDR_WIDTH = 10;
parameter DATA_WIDTH =  75;

logic [ADDR_WIDTH-1:0] addr_reg;

parameter [0:683][DATA_WIDTH-1:0] ROM = {
    //Wall 1
    -75'd1,
    -75'd1,
    -75'd1,
    -75'd1,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,

    //Wall2
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000011111111111111111111111111111111111111111111111111111,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    75'b111100000000000000000000000000000000000000000000000000000000000000000000000,
    -75'd1,
    -75'd1,
    -75'd1,
    -75'd1,

    //Wall 3
    -75'd1,
    -75'd1,
    -75'd1,
    -75'd1,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    

    //Wall 4
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b111111111111111111111111111111111111111111111111111110000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    75'b000000000000000000000000000000000000000000000000000000000000000000000001111,
    -75'd1,
    -75'd1,
    -75'd1,
    -75'd1
};

assign data = ROM[addr];

endmodule