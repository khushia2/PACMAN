module special_walls_6_rom (
    input [1:0] addr,
    output [90:0] data
);

parameter ADDR_WIDTH = 2;
parameter DATA_WIDTH = 91;

logic [ADDR_WIDTH-1:0] addr_reg;

parameter [0:3][DATA_WIDTH-1:0] ROM = {
    //Top 
    -91'd1,
    -91'd1,
    -91'd1,
    -91'd1
};

assign data = ROM[addr];

endmodule