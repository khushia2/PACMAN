module wall_v_rom (
    input [8:0] addr,
    output [3:0] data
);

parameter ADDR_WIDTH = 9;
parameter DATA_WIDTH =  4;

logic [ADDR_WIDTH-1:0] addr_reg;

parameter [0:395][DATA_WIDTH-1:0] ROM = {
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111,
    4'b1111
};

assign data = ROM[addr];

endmodule